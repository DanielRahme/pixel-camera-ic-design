[aimspice]
[description]
2890
Complete-analog-circuit

.include p18_cmos_models.inc
.include p18_model_card.inc

.subckt PhotoDiode VDD N1_R1C1 
I1_R1C1 VDD N1_R1C1 DC Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends PhotoDiode

.subckt OnePixel EXPOSE ERASE NRE OUT vdd vss

.param L1=1.08U
.param W1=1.08U
.param L2=0.36U
.param W2=5.04U
.param L3=0.36U
.param W3=5.04U
.param L4=0.36U
.param W4=5.04U

XD1 vdd N1 PhotoDiode
MN1 N1 EXPOSE N2 vss NMOS L=L1 W=W1
MN2 N2 ERASE vss vss NMOS L=L2 W=W2
CS N2 vss 3pF
MP3 vss N2 N3 vdd PMOS L=L3 W=W3
MP4 N3 NRE OUT vdd PMOS L=L4 W=W4

.ends OnePixel

.param L5=0.36U
.param W5=5.04U
.param L6=0.36U
.param W6=5.04U

XONEPIXEL11 expose erase nre_r1 out1 1 0 ONEPIXEL 
XONEPIXEL12 expose erase nre_r1 out2 1 0 ONEPIXEL
XONEPIXEL21 expose erase nre_r2 out1 1 0 ONEPIXEL
XONEPIXEL22 expose erase nre_r2 out2 1 0 ONEPIXEL
MC1 out1 out1 1 1 PMOS L=L5 W=W5
MC2 out2 out2 1 1 PMOS L=L6 W=W6
CC1 out1 0 3pF
CC2 out2 0 3pF


* This is a parametrized testbench for your pixel circuit array

* You should at least test your circuit with:
*	- current of 50 pA and exposure time 30 ms
*	- current of 750 pA and exposure time 2 ms

* Instructions
* Connect EXPOSE, ERASE, NRE_R1 and NRE_R2 at the right place
* Run a transient simulation with length 60 ms
* Make sure outputs of pixel circuits to ADC are called OUT1 and OUT2
* Make plots of output voltages to ADC (here called OUT1 and OUT2)
* The voltage across internal capacitor (any pixel) is also of interest (here called OUT_SAMPLED1)
* You should also plot the control signals EXPOSE, NRE_R1, NRE_R2 and ERASE

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 30m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

*.plot V(OUT1) V(OUT2) ! signals going to ADC
.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE)
*.plot V(OUT_SAMPLED1)


[dc]
1
vdd
0
1.8
0.1
[tran]
0.001
60m
0
0.1
0
[ana]
4 1
0
1 1
1 1 -0.5 2
5
v(expose)
v(onepixel11:n2)
v(erase)
v(nre_r1)
v(out1)
[end]
