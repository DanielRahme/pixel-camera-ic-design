[aimspice]
[description]
182
MP3-transistor

.include p18_cmos_models.inc
.include p18_model_card.inc

.param L=1.08U
.param W=2.16U

vds vss N3 dc 1.8
vgs N2 N3 dc 0.9

MP3 vss N2 N3 vdd PMOS L=L W=L
[dc]
1
vds
0
1.8
0.1
[ana]
1 1
0
1 1
1 1 -1.2E-05 -5.69448E-48
1
i(vds)
[end]
