`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.10.2019 15:06:34
// Design Name: 
// Module Name: RE_Control
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RE_Control(
    input Exp_increase,
    input Exp_decrease,
    input Init,
    input Reset,
    input Clk,
    output NRE_1,
    output NRE_2,
    output ADC,
    output Expose,
    output Erase
    );
endmodule
