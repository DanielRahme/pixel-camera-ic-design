`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.10.2019 15:06:34
// Design Name: 
// Module Name: Pixel_Electronics
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Pixel_Electronics(
    input NRE_1,
    input NRE_2,
    input ADC,
    input Expose,
    input Erase,
    output ADC_1_out,
    output ADC_2_out
    );
endmodule
